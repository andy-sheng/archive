library ieee;

--clkʱ��Ƶ��Ϊ50MHz
entity other is
port(
);
end other;

architecture behav of other is
begin



end behav;