library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity counting is
port(
	clk: in std_logic;
	cout: out std_logic_vector(7 downto 0));
end counting;

architecture behav of counting is


begin


end behav;