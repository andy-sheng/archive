library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity led is
port(
	clk: in std_logic;--ʱ���ź�
	cout: out std_logic_vector(7 downto 0));--��յLED�����
end led;

architecture behav of led is
begin



end behav;